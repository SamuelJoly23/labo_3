library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

-- |------+------------+---------------+--------------|
-- | Note | Freq (Hz)  | Start address | Sample count |
-- |------+------------+---------------+--------------|
-- | C    | 130.81     | 0x000         | 0x54         |
-- | C#   | 138.59     | 0x054         | 0x4F         |
-- | D    | 146.83     | 0x0A3         | 0x4B         |
-- | D#   | 155.56     | 0x0EE         | 0x46         |
-- | E    | 164.81     | 0x134         | 0x42         |
-- | F    | 174.61     | 0x176         | 0x3F         |
-- | F#   | 185.0      | 0x1B5         | 0x3B         |
-- | G    | 196.0      | 0x1F0         | 0x38         |
-- | G#   | 207.65     | 0x228         | 0x35         |
-- | A    | 220.0      | 0x25D         | 0x32         |
-- | A#   | 233.08     | 0x28F         | 0x2F         |
-- | B    | 246.94     | 0x2BE         | 0x2C         |
-- | C    | 261.63     | 0x2EA         | 0x2A         |
-- |------+------------+---------------+--------------|

entity ROM_qsin is
  port (
    clk_i    : in  std_logic;
    addr_i   : in  std_logic_vector(11 downto 0);
    sample_o : out std_logic_vector(7 downto 0)
    );

end ROM_qsin;

architecture Behavioral of ROM_qsin is
  type ROM_T is array (0 to 787) of std_logic_vector (7 downto 0);
  constant ROM_cst : ROM_T := (
    X"00",  -- Address 0x000 : 130.81 Hz, 0x54 samples
    X"02",
    X"04",
    X"07",
    X"09",
    X"0B",
    X"0E",
    X"10",
    X"12",
    X"15",
    X"17",
    X"19",
    X"1C",
    X"1E",
    X"20",
    X"23",
    X"25",
    X"27",
    X"29",
    X"2C",
    X"2E",
    X"30",
    X"32",
    X"34",
    X"36",
    X"39",
    X"3B",
    X"3D",
    X"3F",
    X"41",
    X"43",
    X"45",
    X"47",
    X"49",
    X"4B",
    X"4D",
    X"4E",
    X"50",
    X"52",
    X"54",
    X"56",
    X"57",
    X"59",
    X"5B",
    X"5C",
    X"5E",
    X"60",
    X"61",
    X"63",
    X"64",
    X"65",
    X"67",
    X"68",
    X"6A",
    X"6B",
    X"6C",
    X"6D",
    X"6E",
    X"70",
    X"71",
    X"72",
    X"73",
    X"74",
    X"75",
    X"76",
    X"76",
    X"77",
    X"78",
    X"79",
    X"79",
    X"7A",
    X"7B",
    X"7B",
    X"7C",
    X"7C",
    X"7D",
    X"7D",
    X"7D",
    X"7E",
    X"7E",
    X"7E",
    X"7E",
    X"7E",
    X"7E",
    X"00",  -- Address 0x054: 138.59Hz, 0x4F samples
    X"02",
    X"05",
    X"07",
    X"0A",
    X"0C",
    X"0F",
    X"11",
    X"13",
    X"16",
    X"18",
    X"1B",
    X"1D",
    X"20",
    X"22",
    X"25",
    X"27",
    X"29",
    X"2C",
    X"2E",
    X"30",
    X"33",
    X"35",
    X"37",
    X"39",
    X"3C",
    X"3E",
    X"40",
    X"42",
    X"44",
    X"46",
    X"48",
    X"4B",
    X"4D",
    X"4F",
    X"50",
    X"52",
    X"54",
    X"56",
    X"58",
    X"5A",
    X"5B",
    X"5D",
    X"5F",
    X"60",
    X"62",
    X"64",
    X"65",
    X"67",
    X"68",
    X"69",
    X"6B",
    X"6C",
    X"6D",
    X"6F",
    X"70",
    X"71",
    X"72",
    X"73",
    X"74",
    X"75",
    X"76",
    X"77",
    X"78",
    X"79",
    X"79",
    X"7A",
    X"7B",
    X"7B",
    X"7C",
    X"7C",
    X"7D",
    X"7D",
    X"7D",
    X"7E",
    X"7E",
    X"7E",
    X"7E",
    X"7E",
    X"00",  -- Adress 0x0A3: 146.83 Hz, 0x4B samples
    X"02",
    X"05",
    X"07",
    X"0A",
    X"0D",
    X"0F",
    X"12",
    X"15",
    X"17",
    X"1A",
    X"1C",
    X"1F",
    X"22",
    X"24",
    X"27",
    X"29",
    X"2C",
    X"2E",
    X"31",
    X"33",
    X"36",
    X"38",
    X"3A",
    X"3D",
    X"3F",
    X"41",
    X"43",
    X"46",
    X"48",
    X"4A",
    X"4C",
    X"4E",
    X"50",
    X"52",
    X"54",
    X"56",
    X"58",
    X"5A",
    X"5C",
    X"5E",
    X"60",
    X"61",
    X"63",
    X"65",
    X"66",
    X"68",
    X"69",
    X"6B",
    X"6C",
    X"6D",
    X"6F",
    X"70",
    X"71",
    X"72",
    X"73",
    X"75",
    X"76",
    X"76",
    X"77",
    X"78",
    X"79",
    X"7A",
    X"7A",
    X"7B",
    X"7C",
    X"7C",
    X"7D",
    X"7D",
    X"7D",
    X"7E",
    X"7E",
    X"7E",
    X"7E",
    X"7E",
    X"00",  -- Address 0x0EE: 155.56Hz, 0x46 samples
    X"02",
    X"05",
    X"08",
    X"0B",
    X"0E",
    X"10",
    X"13",
    X"16",
    X"19",
    X"1B",
    X"1E",
    X"21",
    X"24",
    X"26",
    X"29",
    X"2C",
    X"2E",
    X"31",
    X"33",
    X"36",
    X"38",
    X"3B",
    X"3D",
    X"40",
    X"42",
    X"45",
    X"47",
    X"49",
    X"4C",
    X"4E",
    X"50",
    X"52",
    X"54",
    X"56",
    X"58",
    X"5A",
    X"5C",
    X"5E",
    X"60",
    X"62",
    X"64",
    X"65",
    X"67",
    X"69",
    X"6A",
    X"6C",
    X"6D",
    X"6F",
    X"70",
    X"71",
    X"72",
    X"74",
    X"75",
    X"76",
    X"77",
    X"78",
    X"79",
    X"79",
    X"7A",
    X"7B",
    X"7B",
    X"7C",
    X"7D",
    X"7D",
    X"7D",
    X"7E",
    X"7E",
    X"7E",
    X"7E",
    X"00",  -- Address 0x134: 164.81Hz, 0x42 samples
    X"02",
    X"05",
    X"08",
    X"0B",
    X"0E",
    X"11",
    X"14",
    X"17",
    X"1A",
    X"1D",
    X"20",
    X"23",
    X"26",
    X"29",
    X"2B",
    X"2E",
    X"31",
    X"34",
    X"36",
    X"39",
    X"3C",
    X"3E",
    X"41",
    X"43",
    X"46",
    X"48",
    X"4B",
    X"4D",
    X"4F",
    X"52",
    X"54",
    X"56",
    X"58",
    X"5A",
    X"5D",
    X"5F",
    X"60",
    X"62",
    X"64",
    X"66",
    X"68",
    X"69",
    X"6B",
    X"6D",
    X"6E",
    X"70",
    X"71",
    X"72",
    X"73",
    X"75",
    X"76",
    X"77",
    X"78",
    X"79",
    X"7A",
    X"7A",
    X"7B",
    X"7C",
    X"7C",
    X"7D",
    X"7D",
    X"7E",
    X"7E",
    X"7E",
    X"7E",
    X"00",  -- Address 0x176: 174.61Hz, 0x3F samples
    X"03",
    X"06",
    X"09",
    X"0C",
    X"0F",
    X"12",
    X"16",
    X"19",
    X"1C",
    X"1F",
    X"22",
    X"25",
    X"28",
    X"2B",
    X"2E",
    X"31",
    X"34",
    X"36",
    X"39",
    X"3C",
    X"3F",
    X"42",
    X"44",
    X"47",
    X"49",
    X"4C",
    X"4F",
    X"51",
    X"53",
    X"56",
    X"58",
    X"5A",
    X"5C",
    X"5F",
    X"61",
    X"63",
    X"65",
    X"66",
    X"68",
    X"6A",
    X"6C",
    X"6D",
    X"6F",
    X"70",
    X"72",
    X"73",
    X"74",
    X"76",
    X"77",
    X"78",
    X"79",
    X"7A",
    X"7A",
    X"7B",
    X"7C",
    X"7D",
    X"7D",
    X"7D",
    X"7E",
    X"7E",
    X"7E",
    X"7E",
    X"00",                              -- Adress 0x1B5: 185.0Hz, 0x3B samples
    X"03",
    X"06",
    X"0A",
    X"0D",
    X"10",
    X"14",
    X"17",
    X"1A",
    X"1D",
    X"21",
    X"24",
    X"27",
    X"2A",
    X"2D",
    X"30",
    X"33",
    X"37",
    X"3A",
    X"3C",
    X"3F",
    X"42",
    X"45",
    X"48",
    X"4B",
    X"4D",
    X"50",
    X"52",
    X"55",
    X"57",
    X"5A",
    X"5C",
    X"5E",
    X"61",
    X"63",
    X"65",
    X"67",
    X"69",
    X"6A",
    X"6C",
    X"6E",
    X"70",
    X"71",
    X"73",
    X"74",
    X"75",
    X"76",
    X"78",
    X"79",
    X"7A",
    X"7A",
    X"7B",
    X"7C",
    X"7D",
    X"7D",
    X"7E",
    X"7E",
    X"7E",
    X"7E",
    X"00",                              -- Address 0x1F0: 196.0Hz, 0x38 samples
    X"03",
    X"07",
    X"0A",
    X"0E",
    X"11",
    X"15",
    X"18",
    X"1C",
    X"1F",
    X"23",
    X"26",
    X"29",
    X"2D",
    X"30",
    X"33",
    X"36",
    X"3A",
    X"3D",
    X"40",
    X"43",
    X"46",
    X"49",
    X"4C",
    X"4E",
    X"51",
    X"54",
    X"56",
    X"59",
    X"5B",
    X"5E",
    X"60",
    X"62",
    X"65",
    X"67",
    X"69",
    X"6B",
    X"6D",
    X"6E",
    X"70",
    X"72",
    X"73",
    X"75",
    X"76",
    X"77",
    X"78",
    X"79",
    X"7A",
    X"7B",
    X"7C",
    X"7D",
    X"7D",
    X"7E",
    X"7E",
    X"7E",
    X"7E",
    X"00",  -- Address 0x228: 207.65Hz, 0x35 samples
    X"03",
    X"07",
    X"0B",
    X"0E",
    X"12",
    X"16",
    X"1A",
    X"1D",
    X"21",
    X"25",
    X"28",
    X"2C",
    X"2F",
    X"33",
    X"36",
    X"39",
    X"3D",
    X"40",
    X"43",
    X"46",
    X"49",
    X"4C",
    X"4F",
    X"52",
    X"55",
    X"58",
    X"5A",
    X"5D",
    X"60",
    X"62",
    X"64",
    X"67",
    X"69",
    X"6B",
    X"6D",
    X"6F",
    X"70",
    X"72",
    X"74",
    X"75",
    X"76",
    X"78",
    X"79",
    X"7A",
    X"7B",
    X"7C",
    X"7C",
    X"7D",
    X"7E",
    X"7E",
    X"7E",
    X"7E",
    X"00",                              -- Address 0x25D: 220.0Hz, 0x32 samples
    X"03",
    X"07",
    X"0B",
    X"0F",
    X"13",
    X"17",
    X"1B",
    X"1F",
    X"23",
    X"27",
    X"2A",
    X"2E",
    X"32",
    X"35",
    X"39",
    X"3D",
    X"40",
    X"43",
    X"47",
    X"4A",
    X"4D",
    X"50",
    X"53",
    X"56",
    X"59",
    X"5C",
    X"5F",
    X"61",
    X"64",
    X"66",
    X"68",
    X"6B",
    X"6D",
    X"6F",
    X"71",
    X"72",
    X"74",
    X"75",
    X"77",
    X"78",
    X"79",
    X"7A",
    X"7B",
    X"7C",
    X"7D",
    X"7D",
    X"7E",
    X"7E",
    X"7E",
    X"00",  -- Address 0x28F: 233.08Hz, 0x2F samples
    X"04",
    X"08",
    X"0C",
    X"10",
    X"14",
    X"19",
    X"1D",
    X"21",
    X"25",
    X"29",
    X"2D",
    X"31",
    X"35",
    X"38",
    X"3C",
    X"40",
    X"43",
    X"47",
    X"4A",
    X"4E",
    X"51",
    X"54",
    X"57",
    X"5A",
    X"5D",
    X"60",
    X"63",
    X"65",
    X"68",
    X"6A",
    X"6C",
    X"6E",
    X"70",
    X"72",
    X"74",
    X"76",
    X"77",
    X"78",
    X"7A",
    X"7B",
    X"7C",
    X"7D",
    X"7D",
    X"7E",
    X"7E",
    X"7E",
    X"00",                              -- Address 0x2BE: 246.94, 0x2C samples
    X"04",
    X"08",
    X"0D",
    X"11",
    X"16",
    X"1A",
    X"1E",
    X"23",
    X"27",
    X"2B",
    X"2F",
    X"34",
    X"38",
    X"3C",
    X"3F",
    X"43",
    X"47",
    X"4B",
    X"4E",
    X"52",
    X"55",
    X"58",
    X"5B",
    X"5E",
    X"61",
    X"64",
    X"67",
    X"69",
    X"6C",
    X"6E",
    X"70",
    X"72",
    X"74",
    X"76",
    X"77",
    X"79",
    X"7A",
    X"7B",
    X"7C",
    X"7D",
    X"7D",
    X"7E",
    X"7E",
    X"00",  -- Address 0x2EA: 261.63Hz, 0x2A samples
    X"04",
    X"09",
    X"0E",
    X"12",
    X"17",
    X"1C",
    X"20",
    X"25",
    X"29",
    X"2E",
    X"32",
    X"36",
    X"3B",
    X"3F",
    X"43",
    X"47",
    X"4B",
    X"4E",
    X"52",
    X"56",
    X"59",
    X"5C",
    X"60",
    X"63",
    X"65",
    X"68",
    X"6B",
    X"6D",
    X"70",
    X"72",
    X"74",
    X"76",
    X"77",
    X"79",
    X"7A",
    X"7B",
    X"7C",
    X"7D",
    X"7E",
    X"7E",
    X"7E"
    );

begin

  p_sync : process (clk_i)
  begin
    if rising_edge(clk_i) then
      sample_o <= ROM_cst (to_integer (unsigned (addr_i)));
    end if;
  end process;

end Behavioral;
